--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   12:54:40 04/11/2025
-- Design Name:   
-- Module Name:   /home/student/Desktop/13000123012/ALU/alu_test.vhd
-- Project Name:  ALU
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: alu_rtl
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY alu_test IS
END alu_test;
 
ARCHITECTURE behavior OF alu_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT alu_rtl
    PORT(
         a : IN  std_logic_vector(3 downto 0);
         b : IN  std_logic_vector(3 downto 0);
         s : IN  std_logic_vector(2 downto 0);
         o : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic_vector(3 downto 0) := (others => '0');
   signal b : std_logic_vector(3 downto 0) := (others => '0');
   signal s : std_logic_vector(2 downto 0) := (others => '0');

 	--Outputs
   signal o : std_logic_vector(3 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 

 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: alu_rtl PORT MAP (
          a => a,
          b => b,
          s => s,
          o => o
        );

   -- Clock process definitions


   -- Stimulus process
   stim_proc: process
   begin		
      a<="0010";
		b<="0100";
		s<="000";
		wait for 1 ps;
		a<="0110";
		b<="0100";
		s<="001";
		wait for 1 ps;
		a<="0010";
		b<="0000";
		s<="010";
		wait for 1 ps;
		a<="0110";
		b<="0011";
		s<="011";
		wait for 1 ps;
		a<="0011";
		b<="0100";
		s<="100";
		wait for 1 ps;
		a<="0111";
		b<="0001";
		s<="101";
		wait for 1 ps;
		a<="0011";
		b<="0000";
		s<="110";
		wait for 1 ps;
		a<="0101";
		b<="0011";
		s<="111";
		wait for 1 ps;
   end process;

END;
